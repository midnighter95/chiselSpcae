module And(
  input  a,
         b,
  output z
);

  assign z = a & b;
endmodule
